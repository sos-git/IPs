
module CDK_R512x16(ADDRESS, ROM_OUT, CLOCK, ENABLE);
  input [8:0] ADDRESS;
  input CLOCK, ENABLE;
  output [15:0] ROM_OUT;

endmodule
